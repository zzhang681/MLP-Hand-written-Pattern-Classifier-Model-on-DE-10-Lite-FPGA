
module obs(
	input [31:0] wh1,
	input [31:0] wh2,
	input [31:0] wh3,
	input [31:0] wh4,
	input [31:0] rh1,
	input [31:0] rh2,
	input [31:0] rh3,
	input [31:0] rh4,
	input [31:0] wo1,
	input [31:0] wo2,
	input [31:0] ro1,
	input [31:0] ro2
);



endmodule
